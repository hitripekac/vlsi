arhitecture bla of;
ksdhfdkjshfas
asdfkjhasdfkjhdasf
kjahsfkjdhasf
dsadasda